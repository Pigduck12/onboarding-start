module spi_peripheral (
  
);
